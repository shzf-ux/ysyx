module ysyx_25030085_branch (





);
case(func3)
            3'b000:begin//beq
           
            end
            3'b001:begin//bne
            end
            3'b100:begin//blt
                
            end
            3'b101:begin//bge
                
            end
            3'b110:begin//bltu
                
            end
            3'b111:begin//bgeu
                
            end
            default:begin
                
            end


            endcase   
endmodule
